module camera_module ( 
output reg camera_active 
); 
initial begin camera_active = 1;  
end  
endmodule
